`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: ZJU
// Engineer: tangyi

////////////////////////////////////////////////////////////////////////////////

module PipelineCPU_tb_v;
	// Inputs
	reg clk;
	reg reset;
	// Outputs
	wire [2:0] JumpFlag;
	wire [31:0] Instruction_id;
	wire [31:0] ALU_A;
	wire [31:0] ALU_B;
	wire [31:0] ALUResult;
	wire [31:0] PC;
	wire [31:0] MemDout_mem;
	wire Stall;
	

	// Instantiate the Unit Under Test (UUT)
	PipelineCPU uut (
		.clk(clk), 
		.reset(reset), 
		.JumpFlag(JumpFlag), 
		.Instruction_id(Instruction_id), 
		.ALU_A(ALU_A), 
		.ALU_B(ALU_B), 
		.ALUResult(ALUResult), 
		.PC(PC), 
		.MemDout_mem(MemDout_mem), 
		.Stall(Stall) 
		
	);
      glbl glbl();
	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 0;
        #51     reset = 1;	
                // Wait 100 ns for global reset to finish
	#100 reset=0;
     	#2500 $stop;
	end
	
	always #50 clk=~clk;
      
endmodule

